��- - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 - -  
 - -       F i l e N a m e :                   s p i _ m a s t e r . v h d  
 - -       D e p e n d e n c i e s :           n o n e  
 - -       D e s i g n   S o f t w a r e :     Q u a r t u s   I I   V e r s i o n   9 . 0   B u i l d   1 3 2   S J   F u l l   V e r s i o n  
 - -  
 - -       H D L   C O D E   I S   P R O V I D E D   " A S   I S . "     D I G I - K E Y   E X P R E S S L Y   D I S C L A I M S   A N Y  
 - -       W A R R A N T Y   O F   A N Y   K I N D ,   W H E T H E R   E X P R E S S   O R   I M P L I E D ,   I N C L U D I N G   B U T   N O T  
 - -       L I M I T E D   T O ,   T H E   I M P L I E D   W A R R A N T I E S   O F   M E R C H A N T A B I L I T Y ,   F I T N E S S   F O R   A  
 - -       P A R T I C U L A R   P U R P O S E ,   O R   N O N - I N F R I N G E M E N T .   I N   N O   E V E N T   S H A L L   D I G I - K E Y  
 - -       B E   L I A B L E   F O R   A N Y   I N C I D E N T A L ,   S P E C I A L ,   I N D I R E C T   O R   C O N S E Q U E N T I A L  
 - -       D A M A G E S ,   L O S T   P R O F I T S   O R   L O S T   D A T A ,   H A R M   T O   Y O U R   E Q U I P M E N T ,   C O S T   O F  
 - -       P R O C U R E M E N T   O F   S U B S T I T U T E   G O O D S ,   T E C H N O L O G Y   O R   S E R V I C E S ,   A N Y   C L A I M S  
 - -       B Y   T H I R D   P A R T I E S   ( I N C L U D I N G   B U T   N O T   L I M I T E D   T O   A N Y   D E F E N S E   T H E R E O F ) ,  
 - -       A N Y   C L A I M S   F O R   I N D E M N I T Y   O R   C O N T R I B U T I O N ,   O R   O T H E R   S I M I L A R   C O S T S .  
 - -  
 - -       V e r s i o n   H i s t o r y  
 - -       V e r s i o n   1 . 0   7 / 2 3 / 2 0 1 0   S c o t t   L a r s o n  
 - -           I n i t i a l   P u b l i c   R e l e a s e  
 - -          
 - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
  
 L I B R A R Y   i e e e ;  
 U S E   i e e e . s t d _ l o g i c _ 1 1 6 4 . a l l ;  
 U S E   i e e e . s t d _ l o g i c _ a r i t h . a l l ;  
 U S E   i e e e . s t d _ l o g i c _ u n s i g n e d . a l l ;  
  
 E N T I T Y   s p i _ m a s t e r   I S  
     G E N E R I C (  
         s l a v e s     :   I N T E G E R   : =   8 ;     - - n u m b e r   o f   s p i   s l a v e s  
         d _ w i d t h   :   I N T E G E R   : =   8 ) ;   - - d a t a   b u s   w i d t h  
     P O R T (  
         c l o c k       :   I N           S T D _ L O G I C ;                                                           - - s y s t e m   c l o c k  
         r e s e t _ n   :   I N           S T D _ L O G I C ;                                                           - - a s y n c h r o n o u s   r e s e t  
         e n a b l e     :   I N           S T D _ L O G I C ;                                                           - - i n i t i a t e   t r a n s a c t i o n  
         c p o l         :   I N           S T D _ L O G I C ;                                                           - - s p i   c l o c k   p o l a r i t y  
         c p h a         :   I N           S T D _ L O G I C ;                                                           - - s p i   c l o c k   p h a s e  
         c o n t         :   I N           S T D _ L O G I C ;                                                           - - c o n t i n u o u s   m o d e   c o m m a n d  
         c l k _ d i v   :   I N           I N T E G E R ;                                                               - - s y s t e m   c l o c k   c y c l e s   p e r   1 / 2   p e r i o d   o f   s c l k  
         a d d r         :   I N           I N T E G E R ;                                                               - - a d d r e s s   o f   s l a v e  
         t x _ d a t a   :   I N           S T D _ L O G I C _ V E C T O R ( d _ w i d t h - 1   D O W N T O   0 ) ;     - - d a t a   t o   t r a n s m i t  
         m i s o         :   I N           S T D _ L O G I C ;                                                           - - m a s t e r   i n ,   s l a v e   o u t  
         s c l k         :   B U F F E R   S T D _ L O G I C ;                                                           - - s p i   c l o c k  
         s s _ n         :   B U F F E R   S T D _ L O G I C _ V E C T O R ( s l a v e s - 1   D O W N T O   0 ) ;       - - s l a v e   s e l e c t  
         m o s i         :   O U T         S T D _ L O G I C ;                                                           - - m a s t e r   o u t ,   s l a v e   i n  
         b u s y         :   O U T         S T D _ L O G I C ;                                                           - - b u s y   /   d a t a   r e a d y   s i g n a l  
         r x _ d a t a   :   O U T         S T D _ L O G I C _ V E C T O R ( d _ w i d t h - 1   D O W N T O   0 ) ) ;   - - d a t a   r e c e i v e d  
 E N D   s p i _ m a s t e r ;  
  
 A R C H I T E C T U R E   l o g i c   O F   s p i _ m a s t e r   I S  
     T Y P E   m a c h i n e   I S ( r e a d y ,   e x e c u t e ) ;                                                       - - s t a t e   m a c h i n e   d a t a   t y p e  
     S I G N A L   s t a t e               :   m a c h i n e ;                                                             - - c u r r e n t   s t a t e  
     S I G N A L   s l a v e               :   I N T E G E R ;                                                             - - s l a v e   s e l e c t e d   f o r   c u r r e n t   t r a n s a c t i o n  
     S I G N A L   c l k _ r a t i o       :   I N T E G E R ;                                                             - - c u r r e n t   c l k _ d i v  
     S I G N A L   c o u n t               :   I N T E G E R ;                                                             - - c o u n t e r   t o   t r i g g e r   s c l k   f r o m   s y s t e m   c l o c k  
     S I G N A L   c l k _ t o g g l e s   :   I N T E G E R   R A N G E   0   T O   d _ w i d t h * 2   +   1 ;           - - c o u n t   s p i   c l o c k   t o g g l e s  
     S I G N A L   a s s e r t _ d a t a   :   S T D _ L O G I C ;                                                         - - ' 1 '   i s   t x   s c l k   t o g g l e ,   ' 0 '   i s   r x   s c l k   t o g g l e  
     S I G N A L   c o n t i n u e         :   S T D _ L O G I C ;                                                         - - f l a g   t o   c o n t i n u e   t r a n s a c t i o n  
     S I G N A L   r x _ b u f f e r       :   S T D _ L O G I C _ V E C T O R ( d _ w i d t h - 1   D O W N T O   0 ) ;   - - r e c e i v e   d a t a   b u f f e r  
     S I G N A L   t x _ b u f f e r       :   S T D _ L O G I C _ V E C T O R ( d _ w i d t h - 1   D O W N T O   0 ) ;   - - t r a n s m i t   d a t a   b u f f e r  
     S I G N A L   l a s t _ b i t _ r x   :   I N T E G E R   R A N G E   0   T O   d _ w i d t h * 2 ;                   - - l a s t   r x   d a t a   b i t   l o c a t i o n  
 B E G I N  
     P R O C E S S ( c l o c k ,   r e s e t _ n )  
     B E G I N  
  
         I F ( r e s e t _ n   =   ' 0 ' )   T H E N                 - - r e s e t   s y s t e m  
             b u s y   < =   ' 1 ' ;                                 - - s e t   b u s y   s i g n a l  
             s s _ n   < =   ( O T H E R S   = >   ' 1 ' ) ;         - - d e a s s e r t   a l l   s l a v e   s e l e c t   l i n e s  
             m o s i   < =   ' Z ' ;                                 - - s e t   m a s t e r   o u t   t o   h i g h   i m p e d a n c e  
             r x _ d a t a   < =   ( O T H E R S   = >   ' 0 ' ) ;   - - c l e a r   r e c e i v e   d a t a   p o r t  
             s t a t e   < =   r e a d y ;                           - - g o   t o   r e a d y   s t a t e   w h e n   r e s e t   i s   e x i t e d  
  
         E L S I F ( c l o c k ' E V E N T   A N D   c l o c k   =   ' 1 ' )   T H E N  
             C A S E   s t a t e   I S                               - - s t a t e   m a c h i n e  
  
                 W H E N   r e a d y   = >  
                     b u s y   < =   ' 0 ' ;                           - - c l o c k   o u t   n o t   b u s y   s i g n a l  
                     s s _ n   < =   ( O T H E R S   = >   ' 1 ' ) ;   - - s e t   a l l   s l a v e   s e l e c t   o u t p u t s   h i g h  
                     m o s i   < =   ' Z ' ;                           - - s e t   m o s i   o u t p u t   h i g h   i m p e d a n c e  
                     c o n t i n u e   < =   ' 0 ' ;                   - - c l e a r   c o n t i n u e   f l a g  
  
                     - - u s e r   i n p u t   t o   i n i t i a t e   t r a n s a c t i o n  
                     I F ( e n a b l e   =   ' 1 ' )   T H E N                
                         b u s y   < =   ' 1 ' ;                           - - s e t   b u s y   s i g n a l  
                         I F ( a d d r   <   s l a v e s )   T H E N       - - c h e c k   f o r   v a l i d   s l a v e   a d d r e s s  
                             s l a v e   < =   a d d r ;                   - - c l o c k   i n   c u r r e n t   s l a v e   s e l e c t i o n   i f   v a l i d  
                         E L S E  
                             s l a v e   < =   0 ;                         - - s e t   t o   f i r s t   s l a v e   i f   n o t   v a l i d  
                         E N D   I F ;  
                         I F ( c l k _ d i v   =   0 )   T H E N           - - c h e c k   f o r   v a l i d   s p i   s p e e d  
                             c l k _ r a t i o   < =   1 ;                 - - s e t   t o   m a x i m u m   s p e e d   i f   z e r o  
                             c o u n t   < =   1 ;                         - - i n i t i a t e   s y s t e m - t o - s p i   c l o c k   c o u n t e r  
                         E L S E  
                             c l k _ r a t i o   < =   c l k _ d i v ;     - - s e t   t o   i n p u t   s e l e c t i o n   i f   v a l i d  
                             c o u n t   < =   c l k _ d i v ;             - - i n i t i a t e   s y s t e m - t o - s p i   c l o c k   c o u n t e r  
                         E N D   I F ;  
                         s c l k   < =   c p o l ;                         - - s e t   s p i   c l o c k   p o l a r i t y  
                         a s s e r t _ d a t a   < =   N O T   c p h a ;   - - s e t   s p i   c l o c k   p h a s e  
                         t x _ b u f f e r   < =   t x _ d a t a ;         - - c l o c k   i n   d a t a   f o r   t r a n s m i t   i n t o   b u f f e r  
                         c l k _ t o g g l e s   < =   0 ;                 - - i n i t i a t e   c l o c k   t o g g l e   c o u n t e r  
                         l a s t _ b i t _ r x   < =   d _ w i d t h * 2   +   c o n v _ i n t e g e r ( c p h a )   -   1 ;   - - s e t   l a s t   r x   d a t a   b i t  
                         s t a t e   < =   e x e c u t e ;                 - - p r o c e e d   t o   e x e c u t e   s t a t e  
                     E L S E  
                         s t a t e   < =   r e a d y ;                     - - r e m a i n   i n   r e a d y   s t a t e  
                     E N D   I F ;  
  
                 W H E N   e x e c u t e   = >  
                     b u s y   < =   ' 1 ' ;                 - - s e t   b u s y   s i g n a l  
                     s s _ n ( s l a v e )   < =   ' 0 ' ;   - - s e t   p r o p e r   s l a v e   s e l e c t   o u t p u t  
                      
                     - - s y s t e m   c l o c k   t o   s c l k   r a t i o   i s   m e t  
                     I F ( c o u n t   =   c l k _ r a t i o )   T H E N                  
                         c o u n t   < =   1 ;                                           - - r e s e t   s y s t e m - t o - s p i   c l o c k   c o u n t e r  
                         a s s e r t _ d a t a   < =   N O T   a s s e r t _ d a t a ;   - - s w i t c h   t r a n s m i t / r e c e i v e   i n d i c a t o r  
                         c l k _ t o g g l e s   < =   c l k _ t o g g l e s   +   1 ;   - - i n c r e m e n t   s p i   c l o c k   t o g g l e s   c o u n t e r  
                          
                         - - s p i   c l o c k   t o g g l e   n e e d e d  
                         I F ( c l k _ t o g g l e s   < =   d _ w i d t h * 2   A N D   s s _ n ( s l a v e )   =   ' 0 ' )   T H E N    
                             s c l k   < =   N O T   s c l k ;   - - t o g g l e   s p i   c l o c k  
                         E N D   I F ;  
                          
                         - - r e c e i v e   s p i   c l o c k   t o g g l e  
                         I F ( a s s e r t _ d a t a   =   ' 0 '   A N D   c l k _ t o g g l e s   <   l a s t _ b i t _ r x   +   1   A N D   s s _ n ( s l a v e )   =   ' 0 ' )   T H E N    
                             r x _ b u f f e r   < =   r x _ b u f f e r ( d _ w i d t h - 2   D O W N T O   0 )   &   m i s o ;   - - s h i f t   i n   r e c e i v e d   b i t  
                         E N D   I F ;  
                          
                         - - t r a n s m i t   s p i   c l o c k   t o g g l e  
                         I F ( a s s e r t _ d a t a   =   ' 1 '   A N D   c l k _ t o g g l e s   <   l a s t _ b i t _ r x )   T H E N    
                             m o s i   < =   t x _ b u f f e r ( d _ w i d t h - 1 ) ;                                           - - c l o c k   o u t   d a t a   b i t  
                             t x _ b u f f e r   < =   t x _ b u f f e r ( d _ w i d t h - 2   D O W N T O   0 )   &   ' 0 ' ;   - - s h i f t   d a t a   t r a n s m i t   b u f f e r  
                         E N D   I F ;  
                          
                         - - l a s t   d a t a   r e c e i v e ,   b u t   c o n t i n u e  
                         I F ( c l k _ t o g g l e s   =   l a s t _ b i t _ r x   A N D   c o n t   =   ' 1 ' )   T H E N    
                             t x _ b u f f e r   < =   t x _ d a t a ;                                               - - r e l o a d   t r a n s m i t   b u f f e r  
                             c l k _ t o g g l e s   < =   l a s t _ b i t _ r x   -   d _ w i d t h * 2   +   1 ;   - - r e s e t   s p i   c l o c k   t o g g l e   c o u n t e r  
                             c o n t i n u e   < =   ' 1 ' ;                                                         - - s e t   c o n t i n u e   f l a g  
                         E N D   I F ;  
                          
                         - - n o r m a l   e n d   o f   t r a n s a c t i o n ,   b u t   c o n t i n u e  
                         I F ( c o n t i n u e   =   ' 1 ' )   T H E N      
                             c o n t i n u e   < =   ' 0 ' ;             - - c l e a r   c o n t i n u e   f l a g  
                             b u s y   < =   ' 0 ' ;                     - - c l o c k   o u t   s i g n a l   t h a t   f i r s t   r e c e i v e   d a t a   i s   r e a d y  
                             r x _ d a t a   < =   r x _ b u f f e r ;   - - c l o c k   o u t   r e c e i v e d   d a t a   t o   o u t p u t   p o r t          
                         E N D   I F ;  
                          
                         - - e n d   o f   t r a n s a c t i o n  
                         I F ( ( c l k _ t o g g l e s   =   d _ w i d t h * 2   +   1 )   A N D   c o n t   =   ' 0 ' )   T H E N        
                             b u s y   < =   ' 0 ' ;                           - - c l o c k   o u t   n o t   b u s y   s i g n a l  
                             s s _ n   < =   ( O T H E R S   = >   ' 1 ' ) ;   - - s e t   a l l   s l a v e   s e l e c t s   h i g h  
                             m o s i   < =   ' Z ' ;                           - - s e t   m o s i   o u t p u t   h i g h   i m p e d a n c e  
                             r x _ d a t a   < =   r x _ b u f f e r ;         - - c l o c k   o u t   r e c e i v e d   d a t a   t o   o u t p u t   p o r t  
                             s t a t e   < =   r e a d y ;                     - - r e t u r n   t o   r e a d y   s t a t e  
                         E L S E                                               - - n o t   e n d   o f   t r a n s a c t i o n  
                             s t a t e   < =   e x e c u t e ;                 - - r e m a i n   i n   e x e c u t e   s t a t e  
                         E N D   I F ;  
                      
                     E L S E 	 	 	     - - s y s t e m   c l o c k   t o   s c l k   r a t i o   n o t   m e t  
                         c o u n t   < =   c o u n t   +   1 ;   - - i n c r e m e n t   c o u n t e r  
                         s t a t e   < =   e x e c u t e ;       - - r e m a i n   i n   e x e c u t e   s t a t e  
                     E N D   I F ;  
  
             E N D   C A S E ;  
         E N D   I F ;  
     E N D   P R O C E S S ;    
 E N D   l o g i c ; 